module test (
    output o1,
    output led1,
    input in1
);
    assign o1 = 1'b1;
    assign led1 = in1;
endmodule