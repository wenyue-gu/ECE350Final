module test (
    output o1
);
    assign o1 = 1'b1;

endmodule